LIBRARY IEEE;
LIBRARY ALTERA_MF;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ALTERA_MF.ALTERA_MF_COMPONENTS.ALL;
USE LPM.LPM_COMPONENTS.ALL;

ENTITY UART_OUT_CHK IS

  PORT
  (
	UART_CHK_EN : IN STD_LOGIC;
	NEMPTY		: IN STD_LOGIC;
	IO_DATA		: INOUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END UART_OUT_CHK;

ARCHITECTURE a OF UART_OUT_CHK IS
		
SIGNAL chk_sig		: STD_LOGIC_VECTOR(7 DOWNTO 0);
		
BEGIN
  
  	IO_BUS: LPM_BUSTRI
	GENERIC MAP (
		lpm_width => 8
	)
	PORT MAP (
		data     => chk_sig,
		enabledt => UART_CHK_EN,
		tridata  => IO_DATA
	);
	
	chk_sig <= NEMPTY & NEMPTY & NEMPTY & NEMPTY & NEMPTY & NEMPTY & NEMPTY & NEMPTY;

	
END a;